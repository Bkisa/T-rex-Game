-- author: Furkan Cayci, 2018
-- description: object buffer that holds the objects to display
--    object locations can be controlled from upper level
--    example contains a wall, a rectanble box and a round ball

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity objectbuffer is
    generic (
        OBJECT_SIZE : natural := 16;
        PIXEL_SIZE : natural := 24;
        RES_X : natural := 1280;
        RES_Y : natural := 720
    );
    port (
        video_active       : in  std_logic;
        pixel_x, pixel_y   : in  std_logic_vector(OBJECT_SIZE-1 downto 0);
        object1x, object1y : in  std_logic_vector(OBJECT_SIZE-1 downto 0);
        object2x, object2y : in  std_logic_vector(OBJECT_SIZE-1 downto 0);
        object3x, object3y : in  std_logic_vector(OBJECT_SIZE-1 downto 0);
        object4x, object4y : in  std_logic_vector(OBJECT_SIZE-1 downto 0);
        object5x, object5y : in  std_logic_vector(OBJECT_SIZE-1 downto 0);
        object6x, object6y : in  std_logic_vector(OBJECT_SIZE-1 downto 0);
        object7x, object7y : in  std_logic_vector(OBJECT_SIZE-1 downto 0);
        object8x, object8y : in  std_logic_vector(OBJECT_SIZE-1 downto 0);
        backgrnd_rgb       : in  std_logic_vector(PIXEL_SIZE-1 downto 0);
        rgb                : out std_logic_vector(PIXEL_SIZE-1 downto 0)
    );
end objectbuffer;

architecture rtl of objectbuffer is

    -- x, y coordinates of the trex1
    signal trex_1_x_l : unsigned(OBJECT_SIZE-1 downto 0);
    signal trex_1_x_r : unsigned(OBJECT_SIZE-1 downto 0);
    signal trex_1_y_t : unsigned(OBJECT_SIZE-1 downto 0);
    signal trex_1_y_b : unsigned(OBJECT_SIZE-1 downto 0);

    constant TREX_1 : integer:= 64;

    -- x, y coordinates of the trex2
    signal trex_2_x_l : unsigned(OBJECT_SIZE-1 downto 0);
    signal trex_2_x_r : unsigned(OBJECT_SIZE-1 downto 0);
    signal trex_2_y_t : unsigned(OBJECT_SIZE-1 downto 0);
    signal trex_2_y_b : unsigned(OBJECT_SIZE-1 downto 0);

    constant TREX_2 : integer := 64;
 
    -- x, y coordinates of the trex_dead
    signal trex_dead_x_l : unsigned(OBJECT_SIZE-1 downto 0);
    signal trex_dead_x_r : unsigned(OBJECT_SIZE-1 downto 0);
    signal trex_dead_y_t : unsigned(OBJECT_SIZE-1 downto 0);
    signal trex_dead_y_b : unsigned(OBJECT_SIZE-1 downto 0);

    constant TREX_DEAD : integer :=64;
   
    -- x, y coordinates of the Pterodactyl1
    signal ptero_1_x_l : unsigned(OBJECT_SIZE-1 downto 0);
    signal ptero_1_x_r : unsigned(OBJECT_SIZE-1 downto 0);
    signal ptero_1_y_t : unsigned(OBJECT_SIZE-1 downto 0);
    signal ptero_1_y_b : unsigned(OBJECT_SIZE-1 downto 0);

    constant PTERO_1 : integer :=64;
   
     -- x, y coordinates of the Pterodactyl2
    signal ptero_2_x_l : unsigned(OBJECT_SIZE-1 downto 0);
    signal ptero_2_x_r : unsigned(OBJECT_SIZE-1 downto 0);
    signal ptero_2_y_t : unsigned(OBJECT_SIZE-1 downto 0);
    signal ptero_2_y_b : unsigned(OBJECT_SIZE-1 downto 0);

    constant PTERO_2 : integer :=64;
    
    -- x, y coordinates of the Clouds
    signal cloud_x_l : unsigned(OBJECT_SIZE-1 downto 0);
    signal cloud_x_r : unsigned(OBJECT_SIZE-1 downto 0);
    signal cloud_y_t : unsigned(OBJECT_SIZE-1 downto 0);
    signal cloud_y_b : unsigned(OBJECT_SIZE-1 downto 0);

   	constant CLOUD_SIZE : integer :=64;
  	
   	-- x, y coordinates of the Cactus
   	signal cactus_x_l : unsigned(OBJECT_SIZE-1 downto 0);
   	signal cactus_x_r : unsigned(OBJECT_SIZE-1 downto 0);
   	signal cactus_y_t : unsigned(OBJECT_SIZE-1 downto 0);
   	signal cactus_y_b : unsigned(OBJECT_SIZE-1 downto 0);

   	constant CACTUS_SIZE: integer :=64;

    -- x, y coordinates of the gameover
    signal gameover_x_l : unsigned(OBJECT_SIZE-1 downto 0);
    signal gameover_x_r : unsigned(OBJECT_SIZE-1 downto 0);
    signal gameover_y_t : unsigned(OBJECT_SIZE-1 downto 0);
    signal gameover_y_b : unsigned(OBJECT_SIZE-1 downto 0);

    constant gameover_SIZE: integer :=64;
    
        type rom_type is array (0 to 63) of std_logic_vector(0 to 63);
        
        constant TREX_1_ROM: rom_type :=(
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000011111111111111111111110000000",
            "0000000000000000000000000000000000011111111111111111111110000000",
            "0000000000000000000000000000000011111100111111111111111111110000",
            "0000000000000000000000000000000011111000111111111111111111110000",
            "0000000000000000000000000000000011111000111111111111111111110000",
            "0000000000000000000000000000000011111000111111111111111111110000",
            "0000000000000000000000000000000011111111111111111111111111110000",
            "0000000000000000000000000000000011111111111111111111111111110000",
            "0000000000000000000000000000000011111111111111111111111111110000",
            "0000000000000000000000000000000011111111111111111111111111110000",
            "0000000000000000000000000000000011111111111111111111111111110000",
            "0000000000000000000000000000000011111111111111111111111111110000",
            "0000000000000000000000000000000011111111111111111111111111110000",
            "0000000000000000000000000000000011111111111111111111111111110000",
            "0000000000000000000000000000000011111111111111111111111111110000",
            "0000000000000000000000000000000011111111111111000000000000000000",
            "0000000000000000000000000000000011111111111111000000000000000000",
            "0000000000000000000000000000000011111111111111000000000000000000",
            "0000000000000000000000000000000011111111111111111111100000000000",
            "0000000000000000000000000000000011111111111111111111110000000000",
            "0000000000000000000000000000000011111111111000000000000000000000",
            "0000110000000000000000000000011111111111111000000000000000000000",
            "0000110000000000000000000000011111111111111000000000000000000000",
            "0000110000000000000000000000011111111111111000000000000000000000",
            "0000110000000000000000000111111111111111111000000000000000000000",
            "0000110000000000000000000111111111111111111000000000000000000000",
            "0000111000000000000000000111111111111111111000000000000000000000",
            "0000111110000000000001111111111111111111111111111000000000000000",
            "0000111110000000000001111111111111111111111111111000000000000000",
            "0000111111110000000001111111111111111111111000111000000000000000",
            "0000111111110000000111111111111111111111111000111000000000000000",
            "0000111111110000000111111111111111111111111000111000000000000000",
            "0000111111111000001111111111111111111111111000000000000000000000",
            "0000111111111111111111111111111111111111111000000000000000000000",
            "0000111111111111111111111111111111111111111000000000000000000000",
            "0000111111111111111111111111111111111111111000000000000000000000",
            "0000111111111111111111111111111111111111111000000000000000000000",
            "0000111111111111111111111111111111111111111000000000000000000000",
            "0000001111111111111111111111111111111111111000000000000000000000",
            "0000000111111111111111111111111111111111000000000000000000000000",
            "0000000001111111111111111111111111111111000000000000000000000000",
            "0000000000111111111111111111111111111111000000000000000000000000",
            "0000000000111111111111111111111111111111000000000000000000000000",
            "0000000000000001111111111111111111111000000000000000000000000000",
            "0000000000000001111111111111111111111000000000000000000000000000",
            "0000000000000001111111111111111111111000000000000000000000000000",
            "0000000000000001111111111111111111000000000000000000000000000000",
            "0000000000000001111111111111111111000000000000000000000000000000",
            "0000000000000000111111111111111111000000000000000000000000000000",
            "0000000000000000001111111100011111000000000000000000000000000000",
            "0000000000000000001111111100001111000000000000000000000000000000",
            "0000000000000000001111111000000111000000000000000000000000000000",
            "0000000000000000001111100000000011000000000000000000000000000000",
            "0000000000000000001111100000000011000000000000000000000000000000",
            "0000000000000000001100000000000011111100000000000000000000000000",
            "0000000000000000001100000000000011111100000000000000000000000000",
            "0000000000000000001100000000000000000000000000000000000000000000",
            "0000000000000000001100000000000000000000000000000000000000000000",
            "0000000000000000001111110000000000000000000000000000000000000000",
            "0000000000000000001111110000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000");-- 15
  
               signal trex_1_addr, trex_1_col: unsigned(0 to 5);
               signal trex_1_rom_bit: std_logic;

        constant TREX_2_ROM: rom_type :=(
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000011111111111111111111110000000",
            "0000000000000000000000000000000000011111111111111111111110000000",
            "0000000000000000000000000000000011111100111111111111111111110000",
            "0000000000000000000000000000000011111000111111111111111111110000",
            "0000000000000000000000000000000011111000111111111111111111110000",
            "0000000000000000000000000000000011111000111111111111111111110000",
            "0000000000000000000000000000000011111111111111111111111111110000",
            "0000000000000000000000000000000011111111111111111111111111110000",
            "0000000000000000000000000000000011111111111111111111111111110000",
            "0000000000000000000000000000000011111111111111111111111111110000",
            "0000000000000000000000000000000011111111111111111111111111110000",
            "0000000000000000000000000000000011111111111111111111111111110000",
            "0000000000000000000000000000000011111111111111111111111111110000",
            "0000000000000000000000000000000011111111111111111111111111110000",
            "0000000000000000000000000000000011111111111111111111111111110000",
            "0000000000000000000000000000000011111111111111000000000000000000",
            "0000000000000000000000000000000011111111111111000000000000000000",
            "0000000000000000000000000000000011111111111111000000000000000000",
            "0000000000000000000000000000000011111111111111111111100000000000",
            "0000000000000000000000000000000011111111111111111111110000000000",
            "0000000000000000000000000000000011111111111000000000000000000000",
            "0000110000000000000000000000011111111111111000000000000000000000",
            "0000110000000000000000000000011111111111111000000000000000000000",
            "0000110000000000000000000000011111111111111000000000000000000000",
            "0000110000000000000000000111111111111111111000000000000000000000",
            "0000110000000000000000000111111111111111111000000000000000000000",
            "0000111000000000000000000111111111111111111000000000000000000000",
            "0000111110000000000001111111111111111111111111111000000000000000",
            "0000111110000000000001111111111111111111111111111000000000000000",
            "0000111111110000000001111111111111111111111000111000000000000000",
            "0000111111110000000111111111111111111111111000111000000000000000",
            "0000111111110000000111111111111111111111111000111000000000000000",
            "0000111111111000001111111111111111111111111000000000000000000000",
            "0000111111111111111111111111111111111111111000000000000000000000",
            "0000111111111111111111111111111111111111111000000000000000000000",
            "0000111111111111111111111111111111111111111000000000000000000000",
            "0000111111111111111111111111111111111111111000000000000000000000",
            "0000111111111111111111111111111111111111111000000000000000000000",
            "0000001111111111111111111111111111111111111000000000000000000000",
            "0000000111111111111111111111111111111111000000000000000000000000",
            "0000000001111111111111111111111111111111000000000000000000000000",
            "0000000000111111111111111111111111111111000000000000000000000000",
            "0000000000111111111111111111111111111111000000000000000000000000",
            "0000000000000001111111111111111111111000000000000000000000000000",
            "0000000000000001111111111111111111111000000000000000000000000000",
            "0000000000000001111111111111111111111000000000000000000000000000",
            "0000000000000001111111111111111111000000000000000000000000000000",
            "0000000000000001111111111111111111000000000000000000000000000000",
            "0000000000000000111111111111111111000000000000000000000000000000",
            "0000000000000000001111111100011111000000000000000000000000000000",
            "0000000000000000001111111100011111000000000000000000000000000000",
            "0000000000000000001111110000001111000000000000000000000000000000",
            "0000000000000000001100000000000011000000000000000000000000000000",
            "0000000000000000001100000000000011000000000000000000000000000000",
            "0000000000000000001111110000000011000000000000000000000000000000",
            "0000000000000000001111110000000011000000000000000000000000000000",
            "0000000000000000000000000000000011000000000000000000000000000000",
            "0000000000000000000000000000000011000000000000000000000000000000",
            "0000000000000000000000000000000011111100000000000000000000000000",
            "0000000000000000000000000000000011111100000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000");-- 15

            signal trex_2_addr, trex_2_col: unsigned(0 to 5);
            signal trex_2_rom_bit: std_logic;               

        constant TREX_DEAD_ROM: rom_type :=(
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000111111111111100000000000000000000000000000000000000000000000",
            "0000111111111111100000000000000000000000000000000000000000000000",
            "0000111111111111100000000000000000000000000000000000000000000000",
            "0011111111111111100000000000000000000000000000000000000000000000",
            "0011111111111111100000000000000000000000000000000000000000000000",
            "0011111111111111100000000000000000000000000000000000000000000000",
            "0011111111111111100001000000000000000000000000000000000000000000",
            "0011111111111111100011000000000000000000000000000000000000000000",
            "0011111111111111100011000000000000000000000000000000000000000000",
            "0011111111111111100011000000000000000000000000000000000000000000",
            "0011111111111111100011000000000000000000000000000000000000000000",
            "0011111111111111100011000000011111000000000000000000000000000000",
            "0011111111111111100011000000011111000000000000000000000000000000",
            "0011111111111111100011000000011111000000000000000000000000000000",
            "0011111111111111111111000000011000000000000000000000000000000000",
            "0011111111111111111111000000011000000000000000000000000000000000",
            "0011111111111111111111000000011000000000000000000000000000000000",
            "0011111111111111111111111111111111111111100000000000000000000000",
            "0011111111111111111111111111111111111111100000000000000000000000",
            "0011111111111111111111111111111111111111100000000000000000000000",
            "0011000011111111111111111111111111111111111110000000000000000000",
            "0011000011111111111111111111111111111111111110000000000000000000",
            "0011100011111111111111111111111111111111111110000000000000001100",
            "0011111111111111111111111111111111111111111111110000000000001100",
            "0011111111111111111111111111111111111111111111110000000000001100",
            "0000111111111111111111111111111111111111111111110000000000001100",
            "0000111111111111111111111111111111111111111111111111111111111100",
            "0000111111111111111111111111111111111111111111111111111111111100",
            "0000000000000000000000011111111111111111111111111111110000000000",
            "0000000000000000000000011111111111111111111111111111110000000000",
            "0000000000000000000000011111111111111111111111111111100000000000",
            "0000000000000000000000000011111111111111111111111110000000000000",
            "0000000000000000000000000011111111111111111111111110000000000000",
            "0000000000000000000000000011111111111111111111111110000000000000",
            "0000000000000000000000000011111111111111111111111111100000000000",
            "0000000000000000000000000000011111111111111111111111110000000000",
            "0000000000000000000000000000011111111111111111111111110000001100",
            "0000000000000000000000000000011111111111111111111111111100001100",
            "0000000000000000000000000000011111111111111111111111111100001100",
            "0000000000000000000000000000000011111111111111111111111100001100",
            "0000000000000000000000000000000011111111111111111111111111111100",
            "0000000000000000000000000000000000111111111111111111111111111100",
            "0000000000000000000000000000000000011111111111111110000000000000",
            "0000000000000000000000000000000000011111111111111110000000000000",
            "0000000000000000000000000000000000011111111111111100000000000000",
            "0000000000000000000000000000000000011111111110000000000000000000",
            "0000000000000000000000000000000000011111111110000000000000000000",
            "0000000000000000000000000000000000111111111110000000000000000000",
            "0000000000000000000000000000000111111111111110000000000000000000",
            "0000000000000000000000000000000111111111111110000000000000000000",
            "0000000000000000000000000000000111111111111000000000000000000000",
            "0000000000000000000000000000011111111111110000000000000000000000",
            "0000000000000000000000000000011111111111110000000000000000000000",
            "0000000000000000000000000000111111111111100000000000000000000000",
            "0000000000000000000000011111111111111111000000000000000000000000",
            "0000000000000000000000011111111111111111000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000");-- 15

               signal trex_dead_addr, trex_dead_col: unsigned(0 to 5);
               signal trex_dead_rom_bit: std_logic;
               
        constant CACTUS_ROM: rom_type :=(
            "0000000000000000000000000000111111110000000000000000000000000000",
            "0000000000000000000000000000111111110000000000000000000000000000",
            "0000000000000000000000000000111111110000000000000000000000000000",
            "0000000000000000000000000000111111110000000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000011110000111111111111000011110000000000000000",
            "0000000000000000000011110000111111111111000011110000000000000000",
            "0000000000000000000011110000111111111111000011110000000000000000",
            "0000000000000000000011110000111111111111000011110000000000000000",
            "0000000000000000111111110000111111111111000011110000000000000000",
            "0000000000000000111111110000111111111111000011110000000000000000",
            "0000000000000000111111110000111111111111000011110000000000000000",
            "0000000000000000111111110000111111111111000011110000000000000000",
            "0000000000000000111111110000111111111111000011110000000000000000",
            "0000000000000000111111110000111111111111000011110000000000000000",
            "0000000000000000111111110000111111111111000011110000000000000000",
            "0000000000000000111111110000111111111111000011110000000000000000",
            "0000000000000000111111110000111111111111000011110000000000000000",
            "0000000000000000111111110000111111111111000011110000000000000000",
            "0000000000000000111111110000111111111111000011110000000000000000",
            "0000000000000000111111110000111111111111000011110000000000000000",
            "0000000000000000111111110000111111111111000011110000000000000000",
            "0000000000000000111111110000111111111111000011110000000000000000",
            "0000000000000000111111110000111111111111000011110000000000000000",
            "0000000000000000111111110000111111111111000011110000000000000000",
            "0000000000000000111111111111111111111111111111110000000000000000",
            "0000000000000000111111111111111111111111111111110000000000000000",
            "0000000000000000111111111111111111111111111111110000000000000000",
            "0000000000000000111111111111111111111111111111110000000000000000",
            "0000000000000000000011111111111111111111000000000000000000000000",
            "0000000000000000000011111111111111111111000000000000000000000000",
            "0000000000000000000011111111111111111111000000000000000000000000",
            "0000000000000000000011111111111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000");-- 15
                                 
                 signal cactus_addr, cactus_col: unsigned(0 to 5);
                 signal cactus_rom_bit: std_logic;                 

        constant PTERO_1_ROM: rom_type :=(
            "0000000000000000000000001111111100000000000000000000000000000000",
            "0000000000000000000000001111111100000000000000000000000000000000",
            "0000000000000000000000001111111100000000000000000000000000000000",
            "0000000000000000000000001111111100000000000000000000000000000000",
            "0000000000000000000000001111111111110000000000000000000000000000",
            "0000000000000000000000001111111111110000000000000000000000000000",
            "0000000000000000000000001111111111110000000000000000000000000000",
            "0000000000000000000000001111111111110000000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000000000000000000000111111111111000000000000000000000000",
            "0000000000001111111100000000111111111111111100000000000000000000",
            "0000000000001111111100000000111111111111111100000000000000000000",
            "0000000000001111111100000000111111111111111100000000000000000000",
            "0000000000001111111100000000111111111111111100000000000000000000",
            "0000000011111111111100000000111111111111111111110000000000000000",
            "0000000011111111111100000000111111111111111111110000000000000000",
            "0000000011111111111100000000111111111111111111110000000000000000",
            "0000000011111111111100000000111111111111111111110000000000000000",
            "0000111111111111111100000000111111111111111111111111000000000000",
            "0000111111111111111100000000111111111111111111111111000000000000",
            "0000111111111111111100000000111111111111111111111111000000000000",
            "0000111111111111111100000000111111111111111111111111000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000",
            "1111111111111111111111111111111111111111111111111111000000000000",
            "0000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000000001111111111111111111111111111111100000000",
            "0000000000000000000000001111111111111111111111111111111100000000",
            "0000000000000000000000001111111111111111111111111111111100000000",
            "0000000000000000000000001111111111111111111111111111111100000000",
            "0000000000000000000000000000111111111111111111111111111111110000",
            "0000000000000000000000000000111111111111111111111111111111110000",
            "0000000000000000000000000000111111111111111111111111111111110000",
            "0000000000000000000000000000111111111111111111111111111111110000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000");-- 15
                                 
              signal ptero_1_addr, ptero_1_col: unsigned(0 to 5);
              signal ptero_1_rom_bit: std_logic;                        

        constant PTERO_2_ROM: rom_type :=(
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000001111111100000000000000000000000000000000000000000000",
            "0000000000001111111100000000000000000000000000000000000000000000",
            "0000000000001111111100000000000000000000000000000000000000000000",
            "0000000000001111111100000000000000000000000000000000000000000000",
            "0000000011111111111100000000000000000000000000000000000000000000",
            "0000000011111111111100000000000000000000000000000000000000000000",
            "0000000011111111111100000000000000000000000000000000000000000000",
            "0000000011111111111100000000000000000000000000000000000000000000",
            "0000111111111111111100000000000000000000000000000000000000000000",
            "0000111111111111111100000000000000000000000000000000000000000000",
            "0000111111111111111100000000000000000000000000000000000000000000",
            "0000111111111111111100000000000000000000000000000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000",
            "1111111111111111111111111111111111111111111100000000000000000000",
            "0000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000011111111111111111111111111111111111111111111",
            "0000000000000000000000001111111111111111111111111111111100000000",
            "0000000000000000000000001111111111111111111111111111111100000000",
            "0000000000000000000000001111111111111111111111111111111100000000",
            "0000000000000000000000001111111111111111111111111111111100000000",
            "0000000000000000000000001111111111111111111111111111111111110000",
            "0000000000000000000000001111111111111111111111111111111111110000",
            "0000000000000000000000001111111111111111111111111111111111110000",
            "0000000000000000000000001111111111111111111111111111111111110000",
            "0000000000000000000000001111111111111111111100000000000000000000",
            "0000000000000000000000001111111111111111111100000000000000000000",
            "0000000000000000000000001111111111111111111100000000000000000000",
            "0000000000000000000000001111111111111111111100000000000000000000",
            "0000000000000000000000001111111111110000000000000000000000000000",
            "0000000000000000000000001111111111110000000000000000000000000000",
            "0000000000000000000000001111111111110000000000000000000000000000",
            "0000000000000000000000001111111111110000000000000000000000000000",
            "0000000000000000000000001111111100000000000000000000000000000000",
            "0000000000000000000000001111111100000000000000000000000000000000",
            "0000000000000000000000001111111100000000000000000000000000000000",
            "0000000000000000000000001111111100000000000000000000000000000000",
            "0000000000000000000000001111000000000000000000000000000000000000",
            "0000000000000000000000001111000000000000000000000000000000000000",
            "0000000000000000000000001111000000000000000000000000000000000000",
            "0000000000000000000000001111000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000");-- 15
                                 
             signal ptero_2_addr, ptero_2_col: unsigned(0 to 5);
             signal ptero_2_rom_bit: std_logic;                     

        constant CLOUD_ROM: rom_type :=(
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000001111111111111111111100000000000000000000",
            "0000000000000000000000001111111111111111111100000000000000000000",
            "0000000000000000000000001111111111111111111100000000000000000000",
            "0000000000000000000000001111111111111111111100000000000000000000",
            "0000000000000000000011111111000000000000111111111111111100000000",
            "0000000000000000000011111111000000000000111111111111111100000000",
            "0000000000000000000011111111000000000000111111111111111100000000",
            "0000000000000000000011111111000000000000111111111111111100000000",
            "0000111111111111111111110000000000000000000000000000111111111111",
            "0000111111111111111111110000000000000000000000000000111111111111",
            "0000111111111111111111110000000000000000000000000000111111111111",
            "0000111111111111111111110000000000000000000000000000111111111111",
            "1111111100000000000000000000000000000000000000000000000000001111",
            "1111111100000000000000000000000000000000000000000000000000001111",
            "1111111100000000000000000000000000000000000000000000000000001111",
            "1111111100000000000000000000000000000000000000000000000000001111",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "1111111111111111111111111111111111111111111111111111111111111111",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000");-- 15       

              signal cloud_addr, cloud_col: unsigned(0 to 5);
              signal cloud_rom_bit: std_logic; 
              
        constant gameover : rom_type :=(
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000011111111100000011111000000111000000111001111111111111000",
            "0000000011111111100000011111000000111000001111001111111111111000",
            "0000001111000000000001110011110000111110011111001111000000000000",
            "0000001110000000000001110011110000111110011111001111000000000000",
            "0000011100000000000111000000111000111111111111001111000000000000",
            "0000011100000000000111000000111000111111111111001111000001000000",
            "0000011100001111100111000000111000111111111111001111111111100000",
            "0000011100000111100111111111111000111001101111001111000000000000",
            "0000011100000111100111111111111000111001100111001111000000000000",
            "0000001111000111100111000000111000111000000111001111000000000000",
            "0000001111000111100111000000111000111000000111001111000000000000",
            "0000000011111111100111000000111000111000000111001111111111111000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000001111111110000111000000111000111111111111001111111111100000",
            "0000001111111110000111000000111000111111111111001111111111100000",
            "0000011100000111100111000000111000111000000000001111000001111000",
            "0000011100000111100111000000111000111000000000001111000001111000",
            "0000011100000111100111000000111000111000000000001111000001111000",
            "0000011100000111100111100001111000111100000000001111000001111000",
            "0000011100000111100111110011111000111111111100001111000111111000",
            "0000011100000111100001111111110000111000000000001111111110000000",
            "0000011100000111100001111111110000111000000000001111111110000000",
            "0000011100000111100000011111000000111000000000001111001111100000",
            "0000011100000111100000011111000000111000000000001111001111100000",
            "0000001111111110000000001100000000111111111111001111000111111000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000000000000000000000000000");-- 15
        
                     signal gameover_addr, gameover_col: unsigned(0 to 5);
                     signal gameover_rom_bit: std_logic;
                  
    -- create a 30 pixel vertical wall
    constant WALL_Y_L: integer := 690;
    constant WALL_Y_R: integer := 720;
                  
    -- signals that holds the x, y coordinates
    signal pix_x, pix_y: unsigned (OBJECT_SIZE-1 downto 0);

    signal trex_1_on, trex1, trex_2_on, trex2, trex_dead_on, trexdead, cactus_on, cactuson, cloud_on, cloudon, ptero_1_on, ptero1, ptero_2_on, ptero2, wall_on, gameover_on, gameoveron: std_logic;
    signal trex_1_rgb, trex_2_rgb, trex_dead_rgb, cactus_rgb, cloud_rgb, ptero_1_rgb, ptero_2_rgb, wall_rgb, gameover_rgb: std_logic_vector(23 downto 0);

begin

     pix_x <= unsigned(pixel_x);
     pix_y <= unsigned(pixel_y);
     
     -- draw wall and color
	 wall_on  <= '1' when WALL_Y_L<=pix_y and pix_y<=WALL_Y_R else '0';
	 wall_rgb <= x"FCA207"; -- orange
        
     -- draw trex_1 and color
     trex_1_x_l <= unsigned(object1x);
     trex_1_y_t <= unsigned(object1y);
     trex_1_x_r <= trex_1_x_l + TREX_1 - 1;
     trex_1_y_b <= trex_1_y_t + TREX_1 - 1;
     trex_1_on <= '1' when trex_1_x_l<=pix_x and pix_x<=trex_1_x_r and
                           trex_1_y_t<=pix_y and pix_y<=trex_1_y_b else
                  '0';
     -- trex_1 rgb output
     trex_1_rgb <= x"000000"; -- black
           
     -- draw trex_2 and color
     trex_2_x_l <= unsigned(object2x);
     trex_2_y_t <= unsigned(object2y);
     trex_2_x_r <= trex_2_x_l + TREX_2 - 1;
     trex_2_y_b <= trex_2_y_t + TREX_2 - 1;
     trex_2_on <= '1' when trex_2_x_l<=pix_x and pix_x<=trex_2_x_r and
                           trex_2_y_t<=pix_y and pix_y<=trex_2_y_b else
                 '0';
      -- trex_2 rgb output
     trex_2_rgb <= x"000000"; -- black
            
    -- draw trex_dead and color
     trex_dead_x_l <= unsigned(object3x);
     trex_dead_y_t <= unsigned(object3y);
     trex_dead_x_r <= trex_dead_x_l + TREX_DEAD - 1;
     trex_dead_y_b <= trex_dead_y_t + TREX_DEAD - 1;
     trex_dead_on <= '1' when trex_dead_x_l<=pix_x and pix_x<=trex_dead_x_r and
                              trex_dead_y_t<=pix_y and pix_y<=trex_dead_y_b else
                 '0';
     -- trex_dead rgb output
     trex_dead_rgb <= x"000000"; -- black
    
     -- draw cactus and color
     cactus_x_l <= unsigned(object4x);
     cactus_y_t <= unsigned(object4y);
     cactus_x_r <= cactus_x_l + cactus_SIZE - 1;
     cactus_y_b <= cactus_y_t + cactus_SIZE - 1;
     cactus_on <= '1' when cactus_x_l<=pix_x and pix_x<=cactus_x_r and
                           cactus_y_t<=pix_y and pix_y<=cactus_y_b else
                  '0';
     -- cactus rgb output
     cactus_rgb <= x"00FF00"; -- green
    
     -- draw cloud and color
     cloud_x_l <= unsigned(object5x);
     cloud_y_t <= unsigned(object5y);
     cloud_x_r <= cloud_x_l + cloud_SIZE - 1;
     cloud_y_b <= cloud_y_t + cloud_SIZE - 1;
     cloud_on <= '1' when cloud_x_l<=pix_x and pix_x<=cloud_x_r and
                          cloud_y_t<=pix_y and pix_y<=cloud_y_b else
                 '0';
     -- cloud rgb output
     cloud_rgb <= x"0000FF"; -- blue

     -- draw ptero_1 and color
     ptero_1_x_l <= unsigned(object6x);
     ptero_1_y_t <= unsigned(object6y);
     ptero_1_x_r <= ptero_1_x_l + PTERO_1 - 1;
     ptero_1_y_b <= ptero_1_y_t + PTERO_1- 1;
     ptero_1_on <= '1' when ptero_1_x_l<=pix_x and pix_x<=ptero_1_x_r and
                            ptero_1_y_t<=pix_y and pix_y<=ptero_1_y_b else
                 '0';
     -- ptero_1 rgb output
     ptero_1_rgb <= x"AB00FF"; -- purple
      
     -- draw ptero_2 and color
     ptero_2_x_l <= unsigned(object7x);
     ptero_2_y_t <= unsigned(object7y);
     ptero_2_x_r <= ptero_2_x_l + PTERO_2 - 1;
     ptero_2_y_b <= ptero_2_y_t + PTERO_2 - 1;
     ptero_2_on <= '1' when ptero_2_x_l<=pix_x and pix_x<=ptero_2_x_r and
                            ptero_2_y_t<=pix_y and pix_y<=ptero_2_y_b else
                 '0';
     -- ptero_2 rgb output
     ptero_2_rgb <= x"AB00FF"; -- purple
     
      -- draw gameover and color
     gameover_x_l <= unsigned(object8x);
     gameover_y_t <= unsigned(object8y);
     gameover_x_r <= gameover_x_l + gameover_SIZE - 1;
     gameover_y_b <= gameover_y_t + gameover_SIZE - 1;
     gameover_on <= '1' when gameover_x_l<=pix_x and pix_x<=gameover_x_r and
                            gameover_y_t<=pix_y and pix_y<=gameover_y_b else
                 '0';
     -- gameover rgb output
     gameover_rgb <= x"ff0000"; -- red
     
	 
     -- trex_1 - map current pixel location to ROM addr/col 
     trex_1_addr <= pix_y(5 downto 0) - trex_1_y_t(5 downto 0);
     trex_1_col  <= pix_x(5 downto 0) - trex_1_x_l(5 downto 0);
     trex_1_rom_bit <= TREX_1_ROM(to_integer(trex_1_addr))(to_integer(trex_1_col));
     -- pixel within trex_1
     trex1 <= '1' when trex_1_on='1' and trex_1_rom_bit='1' else '0';
    
     -- trex_2 - map current pixel location to ROM addr/col 
     trex_2_addr <= pix_y(5 downto 0) - trex_2_y_t(5 downto 0);
     trex_2_col  <= pix_x(5 downto 0) - trex_2_x_l(5 downto 0);
     trex_2_rom_bit <= TREX_2_ROM(to_integer(trex_2_addr))(to_integer(trex_2_col));
     -- pixel within trex_2
     trex2 <= '1' when trex_2_on='1' and trex_2_rom_bit='1' else '0';
   
     -- trex_dead - map current pixel location to ROM addr/col 
     trex_dead_addr <= pix_y(5 downto 0) - trex_dead_y_t(5 downto 0);
     trex_dead_col  <= pix_x(5 downto 0) - trex_dead_x_l(5 downto 0);
     trex_dead_rom_bit <= TREX_DEAD_ROM(to_integer(trex_dead_addr))(to_integer(trex_dead_col));
     -- pixel within trex_dead
     trexdead <= '1' when trex_dead_on='1' and trex_dead_rom_bit='1' else '0';     -- !!! trex2 -> trexdead
     
      -- ptero_1 - map current pixel location to ROM addr/col 
     ptero_1_addr <= pix_y(5 downto 0) - ptero_1_y_t(5 downto 0);
     ptero_1_col  <= pix_x(5 downto 0) - ptero_1_x_l(5 downto 0);
     ptero_1_rom_bit <= PTERO_1_ROM(to_integer(ptero_1_addr))(to_integer(ptero_1_col));
     -- pixel within ptero_1
     ptero1 <= '1' when ptero_1_on='1' and ptero_1_rom_bit='1' else '0';
     
    -- ptero_2 - map current pixel location to ROM addr/col 
    ptero_2_addr <= pix_y(5 downto 0) - ptero_2_y_t(5 downto 0);
    ptero_2_col  <= pix_x(5 downto 0) - ptero_2_x_l(5 downto 0);
    ptero_2_rom_bit <= PTERO_2_ROM(to_integer(ptero_2_addr))(to_integer(ptero_2_col));
    -- pixel within ptero_2
    ptero2 <= '1' when ptero_2_on='1' and ptero_2_rom_bit='1' else '0';
   
    -- cloud - map current pixel location to ROM addr/col 
    cloud_addr <= pix_y(5 downto 0) - cloud_y_t(5 downto 0);
    cloud_col  <= pix_x(5 downto 0) - cloud_x_l(5 downto 0);
    cloud_rom_bit <= CLOUD_ROM(to_integer(cloud_addr))(to_integer(cloud_col));
    -- pixel within cloud
    cloudon <= '1' when cloud_on='1' and cloud_rom_bit='1' else '0';
    
    -- cactus - map current pixel location to ROM addr/col 
    cactus_addr <= pix_y(5 downto 0) - cactus_y_t(5 downto 0);
    cactus_col  <= pix_x(5 downto 0) - cactus_x_l(5 downto 0);
    cactus_rom_bit <= CACTUS_ROM(to_integer(cactus_addr))(to_integer(cactus_col));
    -- pixel within cactus
    cactuson <= '1' when cactus_on='1' and cactus_rom_bit='1' else '0';

    -- gameover - map current pixel location to ROM addr/col 
    gameover_addr <= pix_y(5 downto 0) - gameover_y_t(5 downto 0);
    gameover_col  <= pix_x(5 downto 0) - gameover_x_l(5 downto 0);
    gameover_rom_bit <= gameover(to_integer(gameover_addr))(to_integer(gameover_col));
    -- pixel within gameover
    gameoveron <= '1' when gameover_on='1' and gameover_rom_bit='1' else '0';
    
    -- display the image based on who is active
    -- note that the order is important
    process(wall_on,wall_rgb,trex1,trex_1_rgb,trex2,trex_2_rgb,trexdead,trex_dead_rgb,cactuson,cactus_rgb,
	 	    cloudon,cloud_rgb,ptero1,ptero_1_rgb,ptero2,ptero_2_rgb,video_active,backgrnd_rgb, gameoveron, gameover_rgb) is
    begin
		if video_active = '0' then
		  rgb <= x"000000"; --blank
		else
			if trex1='1' then
				rgb <= trex_1_rgb;
			elsif gameoveron='1' then
				rgb <= gameover_rgb; 
			elsif trex2='1' then
				rgb <= trex_2_rgb;   
			elsif trexdead='1' then
				rgb <= trex_dead_rgb;
			elsif cactuson='1' then
				rgb <= cactus_rgb;
			elsif cloudon='1' then
				rgb <= cloud_rgb;   
			elsif ptero1 ='1' then
				rgb <= ptero_1_rgb;
			elsif ptero2='1' then
				rgb <= ptero_2_rgb;
			elsif wall_on='1' then
				rgb <= wall_rgb;         
			else
				rgb <= backgrnd_rgb;
			end if;
	    end if;
   end process;
end rtl;